ruction