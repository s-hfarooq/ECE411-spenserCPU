module reorder_buffer (
    input logic clk,
    input logic rst
);

endmodule : reorder_buffer
