import rv32i_types::*;

module mp4 (
    input clk,
    input rst
);

endmodule : mp4
