module br_pred (
    input logic clk,
    input logic rst
);

endmodule : br_pred
