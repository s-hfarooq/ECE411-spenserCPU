import rv32i_types::*;
import structs::*;
import macros::*;

module cmp_reservation_station (
);

endmodule : cmp_reservation_station
